module EX_MEM (
    input clk,
    input rst,
    
    // info to be passed to MEM
    input [31:0] PC_in,
    input [31:0] inst_in,
    input [4:0] rs1_in,
    input [4:0] rs2_in,
    input [4:0] rd_in,
    input [31:0] alures_in,
    input [31:0] rs2_data_in,
    input Zero_in,

    // corresponding outputs
    output reg[31:0] PC_out,
    output reg[31:0] inst_out,
    output reg[4:0] rs1_out,
    output reg[4:0] rs2_out,
    output reg[4:0] rd_out,
    output reg[31:0] alures_out,
    output reg[31:0] rs2_data_out, 
    output reg Zero_out,
        // the supposed rs2. 
        // when forwarded, this value should be whatever that's passed to alu as rs2.

    // control signals for mem
    input [1:0] MemRead_in,
    output reg[1:0] MemRead_out,
    input [1:0] MemWrite_in,
    output reg[1:0] MemWrite_out,

    // control signals for wb
    input [1:0] RegWrite_in,
    output reg[1:0] RegWrite_out,
    input [1:0] MemtoReg_in,
    output reg[1:0] MemtoReg_out,

    // control for stall
    input stall,
    input flush
);

always @(posedge clk or negedge rst) begin
    if(!rst || flush) 
        begin 
            Zero_out <= 0;
            inst_out <= 0; 
            PC_out <= 0;
            rs1_out <= 0;
            rs2_out <= 0;
            rd_out <= 0;
            alures_out <= 0;
            rs2_data_out <= 0;
            MemRead_out <= 0;
            MemWrite_out <= 0;
            RegWrite_out <= 0;
            MemtoReg_out <= 0; 
        end
    else if(!stall)
        begin
            Zero_out <= Zero_in;
            inst_out <= inst_in; 
            PC_out <= PC_in;
            rs1_out <= rs1_in;
            rs2_out <= rs2_in;
            rd_out <= rd_in;
            rs2_data_out <= rs2_data_in;
            MemRead_out <= MemRead_in;
            MemWrite_out <= MemWrite_in;
            RegWrite_out <= RegWrite_in;
            MemtoReg_out <= MemtoReg_in;
        end

  end

endmodule